`timescale 1ns/1ps

module add_counter_tb;

reg clock;


always @(clock)

BCD7 BCD7
(
    .din        ( din       ),
    .dout       ( dout      )
);

endmodule